magic
tech scmos
timestamp 1638920925
<< nwell >>
rect -22 13 29 32
<< ntransistor >>
rect -2 -11 1 -3
rect 14 -11 17 -3
<< ptransistor >>
rect -2 19 1 26
rect 14 19 17 26
<< ndiffusion >>
rect -5 -11 -2 -3
rect 1 -11 14 -3
rect 17 -11 20 -3
<< pdiffusion >>
rect -4 19 -2 26
rect 1 19 5 26
rect 10 19 14 26
rect 17 19 19 26
<< ndcontact >>
rect -11 -11 -5 -3
rect 20 -11 25 -3
<< pdcontact >>
rect -11 19 -4 26
rect 5 19 10 26
rect 19 19 23 26
<< psubstratepcontact >>
rect -1 -29 4 -22
rect 12 -29 17 -22
<< nsubstratencontact >>
rect -4 39 1 46
rect 10 39 15 46
<< polysilicon >>
rect -2 26 1 38
rect 14 26 17 38
rect -2 -3 1 19
rect 14 -3 17 19
rect -2 -19 1 -11
rect 14 -19 17 -11
<< metal1 >>
rect -11 26 -4 46
rect 1 39 10 46
rect 15 39 31 46
rect 19 26 23 39
rect 5 13 10 19
rect 5 9 25 13
rect 5 8 40 9
rect 20 3 40 8
rect 20 -3 25 3
rect -11 -22 -5 -11
rect -11 -29 -1 -22
rect 4 -29 12 -22
rect 17 -29 31 -22
<< labels >>
rlabel metal1 24 41 24 41 5 vdd
rlabel metal1 23 -26 23 -26 1 gnd
rlabel polysilicon -1 5 -1 5 1 a
rlabel polysilicon 15 -15 15 -15 1 b
rlabel metal1 40 3 40 9 7 y
<< end >>
