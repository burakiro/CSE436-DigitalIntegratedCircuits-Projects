magic
tech scmos
timestamp 1638968460
<< nwell >>
rect -12 6 35 26
<< ntransistor >>
rect -1 -22 1 -16
rect 8 -22 10 -16
rect 18 -22 20 -16
<< ptransistor >>
rect -1 13 1 19
rect 8 13 10 19
rect 18 13 20 19
<< ndiffusion >>
rect -3 -22 -1 -16
rect 1 -22 3 -16
rect 7 -22 8 -16
rect 10 -22 13 -16
rect 17 -22 18 -16
rect 20 -22 25 -16
<< pdiffusion >>
rect -2 13 -1 19
rect 1 13 8 19
rect 10 13 18 19
rect 20 13 25 19
<< ndcontact >>
rect -7 -22 -3 -16
rect 3 -22 7 -16
rect 13 -22 17 -16
rect 25 -22 29 -16
<< pdcontact >>
rect -6 13 -2 19
rect 25 13 29 19
<< polysilicon >>
rect -1 19 1 22
rect 8 19 10 22
rect 18 19 20 22
rect -1 -16 1 13
rect 8 -16 10 13
rect 18 -16 20 13
rect -1 -25 1 -22
rect 8 -25 10 -22
rect 18 -25 20 -22
<< metal1 >>
rect -21 35 49 39
rect -6 19 -2 35
rect 25 -4 29 13
rect 3 -7 41 -4
rect 3 -16 7 -7
rect 25 -16 29 -7
rect -7 -27 -3 -22
rect 13 -27 17 -22
rect -19 -31 51 -27
<< labels >>
rlabel polysilicon 0 -10 0 -10 1 a
rlabel polysilicon 9 -10 9 -10 1 b
rlabel metal1 8 37 8 37 5 vdd
rlabel metal1 5 -29 5 -29 1 gnd
rlabel polysilicon 19 -10 19 -10 1 c
rlabel metal1 41 -7 41 -4 1 y
<< end >>
