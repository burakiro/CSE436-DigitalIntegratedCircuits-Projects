* SPICE3 file created from /home/burakir0/Desktop/hw4/dflip.ext - technology: scmos

.global Vdd Gnd 

.subckt inverter a_n9_n25# a_n14_n6#
M1000 a_n9_n25# a_n14_n6# gnd Gnd nmos w=0.84u l=0.24u
+  ad=0p pd=0u as=0p ps=0u
M1001 a_n9_n25# a_n14_n6# vdd w_n25_10# pmos w=1.68u l=0.24u
+  ad=0p pd=0u as=0p ps=0u
C0 vdd w_n25_10# 0.04fF
C1 a_n9_n25# w_n25_10# 0.05fF
C2 a_n14_n6# w_n25_10# 0.12fF
C3 gnd Gnd 0.18fF
C4 a_n9_n25# Gnd 0.22fF
C5 a_n14_n6# Gnd 0.47fF
C6 vdd Gnd 0.22fF
C7 w_n25_10# Gnd 0.92fF
.ends

.subckt andgate a_n2_n19# gnd a_53_n11# a_14_n51#
M1000 a_1_19# a_n2_n19# vdd w_n22_13# pmos w=0.84u l=0.36u
+  ad=0p pd=0u as=0p ps=0u
M1001 a_53_n11# a_1_19# vdd w_35_12# pmos w=0.84u l=0.6u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_53_n11# a_1_19# gnd Gnd nfet w=0.96u l=0.6u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_1_19# a_14_n51# a_1_n11# Gnd nmos w=0.96u l=0.36u
+  ad=0p pd=0u as=0p ps=0u
M1004 vdd a_14_n51# a_1_19# w_n22_13# pmos w=0.84u l=0.36u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_1_n11# a_n2_n19# gnd Gnd nmos w=0.96u l=0.36u
+  ad=0p pd=0u as=0p ps=0u
C0 gnd a_14_n51# 0.05fF
C1 a_1_19# vdd 0.03fF
C2 a_n2_n19# w_n22_13# 0.15fF
C3 a_1_19# a_14_n51# 0.04fF
C4 w_35_12# vdd 0.06fF
C5 vdd w_n22_13# 0.12fF
C6 a_14_n51# w_n22_13# 0.15fF
C7 w_35_12# a_53_n11# 0.07fF
C8 vdd a_14_n51# 0.05fF
C9 a_1_19# w_35_12# 0.22fF
C10 a_1_19# w_n22_13# 0.07fF
C11 gnd Gnd 0.71fF
C12 a_53_n11# Gnd 0.13fF
C13 a_1_19# Gnd 0.98fF
C14 a_14_n51# Gnd 1.38fF
C15 a_n2_n19# Gnd 0.37fF
C16 vdd Gnd 0.68fF
C17 w_35_12# Gnd 0.63fF
C18 w_n22_13# Gnd 0.87fF
.ends

.subckt nor2gate vdd gnd a_n1_n25# a_1_n22# a_8_n44#
M1000 a_1_13# a_n1_n25# vdd w_n12_6# pmos w=0.72u l=0.24u
+  ad=0p pd=0u as=0p ps=0u
M1001 a_1_n22# a_n1_n25# gnd Gnd nmos w=0.72u l=0.24u
+  ad=0p pd=0u as=0p ps=0u
M1002 gnd a_8_n44# a_1_n22# Gnd nmos w=0.72u l=0.24u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_1_n22# a_8_n44# a_1_13# w_n12_6# pmos w=0.72u l=0.24u
+  ad=0p pd=0u as=0p ps=0u
C0 a_8_n44# a_n1_n25# 0.13fF
C1 a_8_n44# a_1_n22# 0.02fF
C2 w_n12_6# a_n1_n25# 0.11fF
C3 gnd a_8_n44# 0.02fF
C4 w_n12_6# a_1_n22# 0.06fF
C5 a_8_n44# vdd 0.02fF
C6 w_n12_6# vdd 0.06fF
C7 w_n12_6# a_8_n44# 0.15fF
C8 gnd a_1_n22# 0.13fF
C9 gnd Gnd 0.26fF
C10 a_1_n22# Gnd 0.24fF
C11 vdd Gnd 0.46fF
C12 a_8_n44# Gnd 0.78fF
C13 a_n1_n25# Gnd 0.26fF
C14 w_n12_6# Gnd 0.66fF
.ends


* Top level circuit /home/burakir0/Desktop/hw4/dflip

Xinverter_0 a_99_145# d inverter
Xandgate_0 d andgate_0/gnd a_267_n83# clk andgate
Xnor2gate_0 nor2gate_0/vdd nor2gate_0/gnd a_268_159# q q' nor2gate
Xandgate_1 a_99_145# andgate_1/gnd a_268_159# clk andgate
Xnor2gate_1 nor2gate_1/vdd nor2gate_1/gnd a_267_n83# q' q nor2gate
C0 a_267_n83# nor2gate_1/gnd 0.03fF
C1 a_267_n83# q' 0.06fF
C2 andgate_1/gnd a_99_145# 0.09fF
C3 a_268_159# q' 0.00fF
C4 a_268_159# nor2gate_0/gnd 0.03fF
C5 d andgate_0/gnd 0.05fF
C6 a_268_159# q 0.05fF
C7 nor2gate_1/gnd Gnd 0.26fF
C8 q' Gnd 2.87fF
C9 nor2gate_1/vdd Gnd 0.47fF
C10 q Gnd 1.72fF
C11 nor2gate_1/w_n12_6# Gnd 0.66fF 
C12 andgate_1/gnd Gnd 0.71fF
C13 a_268_159# Gnd 1.16fF
C14 andgate_1/a_1_19# Gnd 0.98fF
C15 andgate_1/vdd Gnd 0.68fF 
C16 andgate_1/w_35_12# Gnd 0.63fF 
C17 andgate_1/w_n22_13# Gnd 0.87fF 
C18 nor2gate_0/gnd Gnd 0.26fF
C19 nor2gate_0/vdd Gnd 0.46fF
C20 nor2gate_0/w_n12_6# Gnd 0.66fF 
C21 andgate_0/gnd Gnd 0.71fF
C22 a_267_n83# Gnd 0.96fF
C23 andgate_0/a_1_19# Gnd 0.98fF
C24 clk Gnd 2.98fF
C25 d Gnd 2.36fF
C26 andgate_0/vdd Gnd 0.68fF
C27 andgate_0/w_35_12# Gnd 0.63fF
C28 andgate_0/w_n22_13# Gnd 0.87fF
C29 inverter_0/gnd Gnd 0.18fF
C30 a_99_145# Gnd 1.29fF
C31 inverter_0/vdd Gnd 0.22fF
C32 inverter_0/w_n25_10# Gnd 0.92fF
.end

* INDEPENDANT VOLTAGE SOURCE
*
*Vname +NODE -NODE VALUE
*----- ----- ----- -----
VCC    vdd     0     DC=2.5


* The following two lines are for TRANSIENT analysis
*
*Vname +Node -Node Option T1  V1   T2  V2   T3   V3    T4  V4  T5   V5 
*----- ----- ----- ------ --  --   --  --   ---- --    --  --  ---- -- 
Vina     d     0    PWL(   0   0    4N  0    4.1N 2.5   8N  2.5 8.1N  0  )
Vinb     clk     0    PWL(   0   0    4N  0    4.1N 2.5   8N  2.5 8.1N  0  ) 


*     TSTEP TSTOP
*     ----- -----
.TRAN 0.1N  12N


* The following line is for DC analysis

.DC VIN 0 2.6 0.1


* TEMPERATURE and OPTIONS SETTING

.OPTIONS TEMP=25 reltol = 1e-6 

*MODELS

.include tsmc_cmos025

.END

