* SPICE3 file created from /home/burakir0/Desktop/HW3Integrated/inverter.ext - technology: scmos

M1000 y a gnd Gnd nfet w=0.84u l=0.24u
+  ad=0p pd=0u as=0p ps=0u
M1001 y a vdd w_n25_10# pfet w=1.68u l=0.24u
+  ad=0p pd=0u as=0p ps=0u
C0 y gnd 0.02fF
C1 y w_n25_10# 0.05fF
C2 vdd w_n25_10# 0.04fF
C3 a w_n25_10# 0.12fF
C4 gnd Gnd 0.19fF
C5 y Gnd 0.23fF
C6 a Gnd 0.47fF
C7 vdd Gnd 0.22fF
C8 w_n25_10# Gnd 0.92fF

* INDEPENDANT VOLTAGE SOURCE
*
*Vname +NODE -NODE VALUE
*----- ----- ----- -----
VCC    vdd     0     DC=2.5


* The following two lines are for TRANSIENT analysis
*
*Vname +Node -Node Option T1  V1   T2  V2   T3   V3    T4  V4  T5   V5 
*----- ----- ----- ------ --  --   --  --   ---- --    --  --  ---- -- 
Vina     a     0    PWL(   0   0    4N  0    4.1N 2.5   8N  2.5 8.1N  0  )


*     TSTEP TSTOP
*     ----- -----
.TRAN 0.1N  12N


* The following line is for DC analysis

.DC VIN 0 2.6 0.1


* TEMPERATURE and OPTIONS SETTING

.OPTIONS TEMP=25 reltol = 1e-6 

*MODELS

.include tsmc_cmos025

.END
