magic
tech scmos
timestamp 1635960780
<< nwell >>
rect -22 13 29 32
rect 35 12 70 32
<< ntransistor >>
rect -2 -11 1 -3
rect 14 -11 17 -3
rect 48 -11 53 -3
<< ptransistor >>
rect -2 19 1 26
rect 14 19 17 26
rect 48 19 53 26
<< ndiffusion >>
rect -5 -11 -2 -3
rect 1 -11 14 -3
rect 17 -11 20 -3
rect 41 -11 48 -3
rect 53 -11 58 -3
<< pdiffusion >>
rect -4 19 -2 26
rect 1 19 5 26
rect 10 19 14 26
rect 17 19 19 26
rect 46 19 48 26
rect 53 19 58 26
<< ndcontact >>
rect -11 -11 -5 -3
rect 20 -11 25 -3
rect 35 -11 41 -3
rect 58 -11 64 -3
<< pdcontact >>
rect -11 19 -4 26
rect 5 19 10 26
rect 19 19 23 26
rect 41 19 46 26
rect 58 19 64 26
<< psubstratepcontact >>
rect -1 -29 4 -22
rect 12 -29 17 -22
rect 42 -29 47 -22
rect 56 -29 61 -22
<< nsubstratencontact >>
rect -4 39 1 46
rect 10 39 15 46
rect 44 39 50 46
rect 59 39 65 46
<< polysilicon >>
rect -2 26 1 38
rect 14 26 17 38
rect 48 26 53 38
rect -2 -3 1 19
rect 14 -3 17 19
rect 48 8 53 19
rect 30 4 53 8
rect 48 -3 53 4
rect -2 -19 1 -11
rect 14 -19 17 -11
rect 48 -19 53 -11
<< polycontact >>
rect 25 4 30 8
<< metal1 >>
rect -11 26 -4 46
rect 1 39 10 46
rect 15 39 44 46
rect 50 39 59 46
rect 65 39 70 46
rect 19 26 23 39
rect 41 26 46 39
rect 5 13 10 19
rect 5 8 25 13
rect 20 -3 25 8
rect 58 -3 64 19
rect -11 -22 -5 -11
rect 35 -22 41 -11
rect -11 -29 -1 -22
rect 4 -29 12 -22
rect 17 -29 42 -22
rect 47 -29 56 -22
rect 61 -29 64 -22
<< labels >>
rlabel metal1 24 41 24 41 5 vdd
rlabel metal1 23 -26 23 -26 1 gnd
rlabel polysilicon -1 5 -1 5 1 a
rlabel polysilicon 15 -15 15 -15 1 b
rlabel metal1 59 6 59 6 1 y
<< end >>
