magic
tech scmos
timestamp 1642185088
<< nwell >>
rect -25 10 13 37
<< ntransistor >>
rect -11 -25 -9 -18
<< ptransistor >>
rect -11 17 -9 31
<< ndiffusion >>
rect -17 -21 -11 -18
rect -17 -25 -16 -21
rect -12 -25 -11 -21
rect -9 -22 0 -18
rect -9 -25 4 -22
<< pdiffusion >>
rect -17 29 -11 31
rect -17 25 -16 29
rect -12 25 -11 29
rect -17 17 -11 25
rect -9 24 4 31
rect -9 20 0 24
rect -9 17 4 20
<< ndcontact >>
rect -16 -25 -12 -21
rect 0 -22 4 -18
<< pdcontact >>
rect -16 25 -12 29
rect 0 20 4 24
<< psubstratepcontact >>
rect -16 -37 -12 -30
rect 0 -37 4 -30
<< nsubstratencontact >>
rect -16 39 -12 43
rect 0 39 4 43
<< polysilicon >>
rect -11 31 -9 35
rect -11 -2 -9 17
rect -10 -6 -9 -2
rect -11 -18 -9 -6
rect -11 -28 -9 -25
<< polycontact >>
rect -14 -6 -10 -2
<< metal1 >>
rect -25 39 -16 43
rect -12 39 0 43
rect 4 39 13 43
rect -16 29 -12 39
rect 0 -2 4 20
rect -31 -6 -14 -2
rect 0 -6 12 -2
rect 0 -18 4 -6
rect -16 -30 -12 -25
rect -17 -37 -16 -30
rect -12 -37 0 -30
rect 4 -37 5 -30
<< labels >>
rlabel metal1 -6 -34 -6 -34 1 gnd
rlabel metal1 -6 41 -6 41 5 vdd
<< end >>
