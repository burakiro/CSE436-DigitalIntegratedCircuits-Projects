* SPICE3 file created from andgate.ext - technology: scmos

M1000 a_1_19# a vdd w_n22_13# pmos w=0.84u l=0.36u
+  ad=0p pd=0u as=0p ps=0u
M1001 Y a_1_19# vdd w_35_12# pmos w=0.84u l=0.6u
+  ad=0p pd=0u as=0p ps=0u
M1002 Y a_1_19# 0 0 nmos w=0.96u l=0.6u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_1_19# b a_1_n11# 0 nmos w=0.96u l=0.36u
+  ad=0p pd=0u as=0p ps=0u
M1004 vdd b a_1_19# w_n22_13# pmos w=0.84u l=0.36u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_1_n11# a 0 0 nmos w=0.96u l=0.36u
+  ad=0p pd=0u as=0p ps=0u
C0 w_35_12# a_1_19# 0.22fF
C1 b w_n22_13# 0.15fF
C2 a w_n22_13# 0.15fF
C3 b a_1_19# 0.04fF
C4 w_35_12# vdd 0.06fF
C5 w_35_12# Y 0.07fF
C6 a_1_19# w_n22_13# 0.07fF
C7 vdd w_n22_13# 0.12fF
C8 vdd a_1_19# 0.03fF
C9 0 0 0.71fF
C10 Y 0 0.13fF
C11 a_1_19# 0 0.98fF
C12 b 0 0.37fF
C13 a 0 0.37fF
C14 vdd 0 0.68fF
C15 w_35_12# 0 0.63fF
C16 w_n22_13# 0 0.87fF

* INDEPENDANT VOLTAGE SOURCE
*
*Vname +NODE -NODE VALUE
*----- ----- ----- -----
VCC    vdd     0     DC=2.5


* The following two lines are for TRANSIENT analysis
*
*Vname +Node -Node Option T1  V1   T2  V2   T3   V3    T4  V4  T5   V5 
*----- ----- ----- ------ --  --   --  --   ---- --    --  --  ---- -- 
Vina     a     0    PWL(   0   0    4N  0    4.1N 2.5   8N  2.5 8.1N  0  )
Vinb     b     0    PWL(   0   0    4N  0    4.1N 2.5   8N  2.5 8.1N  0  ) 


*     TSTEP TSTOP
*     ----- -----
.TRAN 0.1N  12N


* The following line is for DC analysis

.DC VIN 0 2.6 0.1


* TEMPERATURE and OPTIONS SETTING

.OPTIONS TEMP=25 reltol = 1e-6 

*MODELS

.include tsmc_cmos025

.END
